module RV32I_X_mem (
    
);
    
endmodule