module ifu_iccm_mem(

)

endmodule
