module RV32I_X (
    
);
    
endmodule