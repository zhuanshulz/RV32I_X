module exe (
    
);
    
endmodule