module dec (
    
);
    
endmodule