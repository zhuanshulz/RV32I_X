module lsu (
    
);
    
endmodule