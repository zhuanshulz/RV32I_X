module dccm_mem(

);

endmodule
