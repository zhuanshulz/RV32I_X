module mem (
    
);
    
endmodule